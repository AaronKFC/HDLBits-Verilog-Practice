module top_module(
    input clk,
    input reset,    // Synchronous reset to OFF
    input j,
    input k,
    output out); //  

    // Solution1 (My implementation) (almost the same as Solution2)
    parameter OFF=0, ON=1;
    reg state, next_s;
    
    always @(*) begin
        case(state)
            OFF: next_s <= j ? ON:OFF;
            ON: next_s <= k ? OFF:ON;
        endcase
    end
    
    always @(posedge clk) begin
        if(reset) state <=OFF;
        else state <= next_s;
    end
    assign out = (state == ON);

    ///////////////////////////////////////////////
    // Solution2
    parameter OFF = 0, ON = 1; 
    reg state, next_state;

    always @(*) begin
        // State transition logic
        case (state)
            ON: next_state <= k ? OFF : ON;
            OFF: next_state <= j ? ON : OFF;
        endcase
    end

    always @(posedge clk) begin
        // State flip-flops with synchronous reset
        if (reset) begin
            state <= OFF;
        end
        else begin
            state <= next_state;
        end
    end

    // Output logic
    // assign out = (state == ...);
    assign out = (state == ON);

endmodule
